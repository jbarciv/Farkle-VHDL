-- Esto es un comentario en VHDL
-- Otro comentario